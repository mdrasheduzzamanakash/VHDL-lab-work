
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity fullAdr is
end fullAdr;

architecture Behavioral of fullAdr is

begin


end Behavioral;

